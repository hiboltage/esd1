
module nios_system (
	clk_clk,
	out_wave_out_wave,
	reset_reset_n);	

	input		clk_clk;
	output		out_wave_out_wave;
	input		reset_reset_n;
endmodule
