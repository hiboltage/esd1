
module nios_system (
	clk_clk,
	key_export,
	leds_export);	

	input		clk_clk;
	input		key_export;
	output	[9:0]	leds_export;
endmodule
